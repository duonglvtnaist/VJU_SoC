`define BITWIDTH        8
`define FULLBITWIDTH    32
`define ADDR_WIDTH      18
`define MODE_ADDR_WIDTH 2


`define AXI_DATA_WIDTH              32